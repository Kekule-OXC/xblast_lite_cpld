-- Code your testbench here
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

-- entity declaration for your testbench.Dont declare any ports here
ENTITY LPCMod_tb IS
END LPCMod_tb;

ARCHITECTURE behavior OF LPCMod_tb IS
   -- Component Declaration for the Unit Under Test (UUT)
    COMPONENT entity_lpcmod is  --'test' is the name of the module needed to be tested.
--just copy and paste the input and output ports of your module as such.
    port (
        pin_xbox_n_lrst : in std_logic;                         -- Xbox-side Reset signal
        pin_xbox_lclk : in std_logic ;                          -- Xbox-side CLK, goes to flash chip too
        pinout4_xbox_lad : inout std_logic_vector(3 downto 0);  -- Xbox-side LPC IO
        pinout4_flash_lad :inout std_logic_vector(3 downto 0);  -- Flash-side LPC IO
        pout_xbox_lframe : out std_logic;                       -- Only goes to tri-state buffer for LFRAME signal control on Xbox motherboard
        pout_flash_lframe : out std_logic;                      -- Only goes to flash chip. Is generated by code logic.
        pout_xbox_d0 : out std_logic ;                          -- D0 control on Xbox motherbord. Useful on all motherboards but 1.6(b) should really USE L1 instead!
        pout_xbox_a19control : out std_logic;                   -- Controls if buffer is tri-stated or driving pout_xbox_a19.
        pout_xbox_a19 : out std_logic;                          -- TSOP bank control. Hooks to Xbox's TSOP pout_xbox_a19.
        pout_xbox_a15 : out std_logic ;                         -- Xbox TSOP pout_xbox_a15 control signal.
        pin_manual_bank1 : in std_logic;                        -- First switch input. Used to split 1MB flash in 2 512KB banks
        pin_manual_bank2 : in std_logic;                        -- Second switch.
        p6out_lcd_data : out std_logic_vector(5 downto 0);      -- Contains R/S, E and D4-D7. R/W is set on W.
        pout_lcd_contrast: out std_logic;                       -- For LCD contrast
        pout_lcd_backlight: out std_logic;                      -- LCD backlight control.
        pout_enable_5v: out std_logic;                          -- Controls onboard +5V switch
        p4out_gpo: out std_logic_vector(3 downto 0);            -- General Purpose Outputs
        p2in_gpi: in std_logic_vector(1 downto 0);              -- General Purpose Inputs
        pout_n_onboard_led : out std_logic                      -- Status led on board
    );
    END COMPONENT entity_lpcmod;
    
    signal pin_xbox_n_lrst : std_logic := '0';
    signal pin_xbox_lclk : std_logic := '0';
    signal pinout4_xbox_lad : std_logic_vector(3 downto 0) := "1111";
    signal pinout4_flash_lad : std_logic_vector(3 downto 0) := "0000";
    signal pout_xbox_lframe : std_logic := '1';
    signal pout_flash_lframe : std_logic;
    signal pout_xbox_d0 : std_logic := '1';
    signal pout_xbox_a19control : std_logic := '1';
    signal pout_xbox_a19 : std_logic := '1';
    signal pout_xbox_a15 : std_logic := '1';
    signal pin_manual_bank1 : std_logic := '1';
    signal pin_manual_bank2 : std_logic := '1';
    signal p6out_lcd_data : std_logic_vector(5 downto 0) := "000000";      --Contains R/S, E and D4-D7. R/W is set on W.
    signal pout_lcd_contrast: std_logic := '0';    --For LCD contrast
    signal pout_lcd_backlight: std_logic:= '0'; --LCD backlight control
    signal pout_enable_5v : std_logic;
    signal p4out_gpo : std_logic_vector(3 downto 0);
    signal p2in_gpi : std_logic_vector(1 downto 0);
    signal pout_n_onboard_led : std_logic;
    
    constant clk_period : time := 30 NS;
    
BEGIN
    -- Instantiate the Unit Under Test (UUT)
   uut: entity_lpcmod PORT MAP (
     pin_xbox_n_lrst,
     pin_xbox_lclk,
     pinout4_xbox_lad,
     pinout4_flash_lad,
     pout_xbox_lframe,
     pout_flash_lframe,
     pout_xbox_d0,
     pout_xbox_a19control,
     pout_xbox_a19,
     pout_xbox_a15,
     pin_manual_bank1,
     pin_manual_bank2
     p6out_lcd_data,
     pout_lcd_contrast,
     pout_lcd_backlight,
     pout_enable_5v,
     p4out_gpo,
     p2in_gpi,
     pout_n_onboard_led
     ); 
        
   -- Clock process definitions( clock with 50% duty cycle is generated here.
   clk_process :process
   begin
        pin_xbox_lclk <= '0';
        wait for clk_period/2;
        pin_xbox_lclk <= '1';
        wait for clk_period/2;
   end process;       
   
   
stim_proc: process
    begin    
        pin_xbox_n_lrst <= '0';
        pin_manual_bank1 <= '1'; -- Default state because of pull-up
        pin_manual_bank2 <= '1'; -- Default state because of pull-up
        pinout4_flash_lad <= "ZZZZ";
        wait for clk_period;        --30 ns delay
        wait for clk_period;
        wait for clk_period;
        wait for 22 NS;         --Arbitrary delay induced on further data stimulation. In reality, the Xbox sets it's data for the next rising edge around 9 NS after the preceding rising edge of said data.
        pin_xbox_n_lrst <= '1';
        wait for clk_period;
        wait for clk_period;
        
        
        
        -- Test LPC mem write
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period; 
        pinout4_flash_lad <= X"F";  --TARA2
        pinout4_xbox_lad <= "ZZZZ";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ";
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0110"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"2";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period; 
        pinout4_flash_lad <= X"F";  --TARA2
        pinout4_xbox_lad <= "ZZZZ";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ";
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        -- Test LPC mem read
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0100"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_flash_lad <= X"F";  --TARA2
        pinout4_xbox_lad <= "ZZZZ";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= x"2";   --DATA1
        wait for clk_period;
        pinout4_flash_lad <= x"5";   --DATA2
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ";  
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0100"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_flash_lad <= X"F";  --TARA2
        pinout4_xbox_lad <= "ZZZZ";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_flash_lad <= x"A";   --DATA2
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ";  
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        -- Test LPC IO write
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC       IO
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr7     LCD
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"3";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;    
        pinout4_xbox_lad <= x"0";   --addr7     LCD
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"6";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;    
        pinout4_xbox_lad <= x"0";   --addr7     LCD
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"5";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"1";   --addr7     Backlight
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"3";   --addr7     Contrast
        wait for clk_period;
        pinout4_xbox_lad <= x"1";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"4";   --addr7     MCU-4
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"2";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"6";   --addr7     MCU-6
        wait for clk_period;
        pinout4_xbox_lad <= x"1";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"6";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"3";   --addr7     Contrast
        wait for clk_period;
        pinout4_xbox_lad <= x"1";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr7     MCU-7
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"A";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        -- Test LPC mem read once more
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0100"; --CYC           Flash read
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr0
        wait for clk_period;
        pinout4_xbox_lad <= "1111"; --addr1
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr2
        wait for clk_period;
        pinout4_xbox_lad <= "0000"; --addr3
        wait for clk_period;
        pinout4_xbox_lad <= x"1";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"2";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"3";   --addr6
        wait for clk_period;
        pinout4_xbox_lad <= x"4";   --addr7
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARA1
        wait for clk_period;
        pinout4_flash_lad <= X"F";  --TARA2
        pinout4_xbox_lad <= "ZZZZ";
        wait for clk_period;
        pinout4_flash_lad <= "0000"; --SYNC
        wait for clk_period;
        pinout4_flash_lad <= x"3";   --DATA1
        wait for clk_period;
        pinout4_flash_lad <= x"4";   --DATA2
        wait for clk_period;
        pinout4_flash_lad <= X"F";   --TARB1
        wait for clk_period;
        pinout4_flash_lad <= "ZZZZ";  
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        
        
        
        -- Test LPC io write once more
        pinout4_xbox_lad <= "0000"; --Start!
        wait for clk_period;
        pinout4_xbox_lad <= "0010"; --CYC
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --addr4
        wait for clk_period;
        pinout4_xbox_lad <= x"7";   --addr5
        wait for clk_period;
        pinout4_xbox_lad <= x"0";   --addr6
        wait for clk_period;    
        pinout4_xbox_lad <= x"0";   --addr7     LCD
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --DATA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F";   --DATA2
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA1
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARA2, stays at 0xF because of pullups
        wait for clk_period;
        --SYNC
        wait for clk_period;
        pinout4_xbox_lad <= x"F"; --TARB1, stays at 0xF because of pullups
        wait for clk_period;
        pinout4_xbox_lad <= X"F";   --TARB2
        wait for clk_period;
        wait for clk_period;
        wait for clk_period;
        ASSERT FALSE REPORT "Test done." SEVERITY NOTE;
        wait;
    end process;

END behavior;
