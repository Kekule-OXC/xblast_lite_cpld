-- Xbox Original modchip code for XBlast-compatible firmware support and extra hw-specific features
-- Copyright (C) 2019  Benjamin Fiset-Deschênes

-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU Lesser General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- any later version.

-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU Lesser General Public License for more details.

-- You should have received a copy of the GNU Lesser General Public License
-- along with this program.  If not, see <https://www.gnu.org/licenses/>.


-- Interface Xbox LPC to SST49LF080A flash device
-- Extra software control for bank switching
-- Support for parallel character LCD with contrast and backlight software control
-- Support for onboard TSOP split software control (Xbox TSOP A19)
-- Support for onboard TSOP recover a la Matrix/Chameleon (Xbox TSOP A15)
-- Support for general purpose input and output pins
-- Support Xodus software control scheme
-- Basic Chihiro MediaBoard spoof
-- Originally designed for XC9572XL CPLD

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;


-- ----------------------------------------
entity entity_lpcmod is
-- ----------------------------------------
    port (
        pin_xbox_n_lrst : in std_logic;                         -- Xbox-side Reset signal
        pin_xbox_lclk : in std_logic ;                          -- Xbox-side CLK, goes to flash chip too
        pinout4_xbox_lad : inout std_logic_vector(3 downto 0);  -- Xbox-side LPC IO
        pinout4_flash_lad :inout std_logic_vector(3 downto 0);  -- Flash-side LPC IO
        pout_xbox_lframe : out std_logic;                       -- Only goes to tri-state buffer for LFRAME signal control on Xbox motherboard
        pout_flash_lframe : out std_logic;                      -- Only goes to flash chip. Is generated by code logic.
        pout_xbox_d0 : out std_logic ;                          -- D0 control on Xbox motherbord. Useful on all motherboards but 1.6(b) should really USE L1 instead!
        pout_xbox_a19control : out std_logic;                   -- Controls if buffer is tri-stated or driving pout_xbox_a19.
        pout_xbox_a19 : out std_logic;                          -- TSOP bank control. Hooks to Xbox's TSOP pout_xbox_a19.
        pout_xbox_a15 : out std_logic ;                         -- Xbox TSOP pout_xbox_a15 control signal.
        pin_manual_bank1 : in std_logic;                        -- First switch input. Used to split 1MB flash in 2 512KB banks
        pin_manual_bank2 : in std_logic;                        -- Second switch.
        p6out_lcd_data : out std_logic_vector(5 downto 0);      -- Contains R/S, E and D4-D7. R/W is set on W.
        pout_lcd_contrast: out std_logic;                       -- For LCD contrast
        pout_lcd_backlight: out std_logic;                      -- LCD backlight control.
        pout_enable_5v: out std_logic;                          -- Controls onboard +5V switch
        p4out_gpo: out std_logic_vector(3 downto 0);            -- General Purpose Outputs
        p2in_gpi: in std_logic_vector(1 downto 0);              -- General Purpose Inputs
        pout_n_onboard_led : out std_logic                      -- Status led on board
    );
end entity_lpcmod;

-- ----------------------------------------
architecture arch_lpcmod of entity_lpcmod is
-- ----------------------------------------
--**+ constants +***
    constant c_FALSE_STD: std_logic := '0';
    constant c_TRUE_STD: std_logic := '1';
    
    constant c_RST_ASSERTED: std_logic := '0';
    
    constant c_LAD_IDLE_PATTERN: std_Logic_vector := "1111";
    constant c_LAD_INPUT_PATTERN: std_Logic_vector := "ZZZZ";

    constant c_LAD_START_PATTERN: std_Logic_vector := "0000";
    constant c_CYC_MEM_PREFIX: std_Logic_vector := "01";
    constant c_CYC_IO_PREFIX: std_Logic_vector := "00";
    
    constant c_CYC_DIRECTION_READ: std_logic := '0';
    constant c_CYC_DIRECTION_WRITE: std_logic := '1';
    
    constant c_LAD_ADDR_PATTERN1: std_Logic_vector := "1111";
    
    constant c_LAD_ST49LF080A_ADDR_PATTERN1: std_Logic_vector := "1110"; -- 1st (highest) addr nibble. Fixed addr bit & MSB Chip ID
    constant c_LAD_ST49LF080A_ADDR_PATTERN2: std_Logic_vector := "0100"; -- 2nd addr nibble. chip ID bit(2) & Memory access signal bit & 2 LSB Chip ID.
    
    constant c_DEV_ID_LOW_NIBBLE: std_logic_vector := "0101";  -- SmartXX OPX/XBlast Lite ID
    constant c_DEV_ID_HIGH_NIBBLE: std_logic_vector := "0001"; -- XBlast gen1
    
    constant c_MEDIABOARD_SPOOF_ID_LOW_NIBBLE: std_logic_vector := "0000";   -- FPGA MediaBoard revision. Change to X"1" to spoof ASIC revision.
    constant c_MEDIABOARD_SPOOF_ID_HIGH_NIBBLE: std_logic_vector := "0000";  -- MediaBoard spoof (very basic...).
    
    constant c_LAD_IOREG_PATTERN1: std_Logic_vector := "1111";
    constant c_LAD_XODUS_PATTERN1: std_Logic_vector := "0000";
    constant c_LAD_MBOARD_PATTERN1: std_Logic_vector := "0100";
    constant c_LAD_IOREG_PATTERN2: std_Logic_vector := "0111";
    constant c_LAD_XODUS_PATTERN2: std_Logic_vector := "0000";
    constant c_LAD_IOREG_PATTERN3: std_Logic_vector := "0000";
    constant c_LAD_XODUS_PATTERN3: std_Logic_vector := "1111";
    
    constant c_LAD_PATTERN_SYNC: std_Logic_vector := "0000";
    
    constant c_FSM_COUNT_RESET: integer := 0;
    constant c_FSM_COUNT_IO_START_OFFSET: integer := 4;
    constant c_FSM_DATA_WRITE_LO_NIBBLE_OFFSET: integer := 0;
    constant c_FSM_DATA_WRITE_HI_NIBBLE_OFFSET: integer := 1;
    
    constant c_FSM_ADDR_SEQ_NIBBLE0: integer := 0;
    constant c_FSM_ADDR_SEQ_NIBBLE1: integer := 1;
    constant c_FSM_ADDR_SEQ_NIBBLE2: integer := 2;
    constant c_FSM_ADDR_SEQ_NIBBLE3: integer := 3;
    constant c_FSM_ADDR_SEQ_NIBBLE4: integer := 4;
    constant c_FSM_ADDR_SEQ_NIBBLE5: integer := 5;
    constant c_FSM_ADDR_SEQ_NIBBLE6: integer := 6;
    constant c_FSM_ADDR_SEQ_NIBBLE7: integer := 7;
    constant c_FSM_ADDR_SEQ_MAX_COUNT: integer := c_FSM_ADDR_SEQ_NIBBLE7;
    constant c_FSM_DATA_SEQ_MAX_COUNT: integer := c_FSM_ADDR_SEQ_NIBBLE6;
    
    constant c_LAD_IOREG_RD_DEV_ID: std_Logic_vector := X"1";
    constant c_LAD_IOREG_RD_MEDIABOARD_RAM: std_Logic_vector := X"4";   -- MediaBoard DIMM size spoof
    constant c_LAD_IOREG_RD_IO: std_Logic_vector := X"D";
    constant c_LAD_IOREG_RD_XODUSID: std_Logic_vector := X"E";
    constant c_LAD_IOREG_RD_STATUS: std_Logic_vector := X"F";
    constant c_LAD_IOREG_RD_MEDIABOARD_ID: std_Logic_vector := X"F";
    constant c_LAD_IOREG_MEDIABOARD_SPOOF_GENERIC: std_Logic_vector := X"C";
    
    constant c_LAD_IOREG_WR_LCD_DATA: std_Logic_vector := X"0";
    constant c_LAD_IOREG_WR_LCD_BACKLIGHT: std_Logic_vector := X"1";
    constant c_LAD_IOREG_WR_LCD_CONTRAST: std_Logic_vector := X"3";
    constant c_LAD_IOREG_WR_OUTPUTS: std_Logic_vector := X"D";
    constant c_LAD_IOREG_WR_CTRL: std_Logic_vector := X"F";
    
    constant c_FSM_DATA_SEQ_TARA2_READ: integer := 1;
    constant c_FSM_DATA_SEQ_TARA2_WRITE: integer := 3;

    constant c_FSM_DATA_SEQ_DATA1_READ: integer := 3;
    constant c_FSM_DATA_SEQ_DATA2_READ: integer := 4;
    
    constant c_FSM_DATA_SEQ_SYNC_READ: integer := 2;
    constant c_FSM_DATA_SEQ_SYNC_WRITE: integer := 4;
    
    constant c_GPO_RESET: std_Logic_vector := "0000";
    
    constant c_LCD_REG_DATA_RESET: std_Logic_vector := "000";
    
    constant c_MEDIABOARD_SPOOF_RAM_SIZE: std_Logic_vector := X"3";   -- MediaBoard DIMM size 1024MB
    
    constant c_PWM_COUNTER_RESET_VALUE: std_Logic_vector := "000000";
    constant c_PWM_COUNTER_MAX_VALUE: std_Logic_vector := "111111";
    constant c_NULL_DUTY_CYCLE: std_Logic_vector := "000000";
    
    constant c_BANK_CTRL_OS_BANK: std_Logic_vector := "11";

--***+ types
    -- Regroup the necessary 17 cycle for a single byte of data transfer (both in R/W).
    type LPC_FSM is (
        LPC_FSM_WAIT_START,  -- 0000 read, occurs with LFRAME output asserted. Active while idle and on START frame (1/17 cycle)
        LPC_FSM_GET_CYC,     -- next nibble is CYCTYPE, only interested in 010x (mem rd) and 011x (mem write), size is always 1 byte for memory. Active 1/17 cycle.
        LPC_FSM_GET_ADDR,    -- 8 nibbles of address, most significant nibble first. Active 8/17 cycles
        LPC_FSM_DATA         -- TAR,SYNC and DATA transfer sequences. Active 7/17 cycles.
    );                       -- For a total of 17 cycles :)


--***+ signals
    signal s_fsm_counter : integer range c_FSM_COUNT_RESET to c_FSM_ADDR_SEQ_MAX_COUNT; -- Used for addresses resolution and LPC_FSM_DATA state counter.
    signal s_lpc_fsm_state : LPC_FSM := LPC_FSM_WAIT_START;                             --2 bit state descriptor, unless you add entries to "LPC_FSM".
    signal s_lad_dir : std_logic;                                                       -- 0 for Flash to Xbox(LPC read)
    signal s_io_cyc : boolean;
    signal s_lframe : std_logic;                                                        -- Internal signal to control pout_flash_lframe and pout_xbox_lframe at the same time.
    signal s6_duty_cycle_backlight : std_Logic_vector(5 downto 0) := c_NULL_DUTY_CYCLE; 
    signal s6_duty_cycle_contrast : std_Logic_vector(5 downto 0) := c_NULL_DUTY_CYCLE;
    signal s6_pwm_counter : std_logic_vector(5 downto 0) := c_PWM_COUNTER_RESET_VALUE;
    signal s4_io_reg_addr : std_logic_vector(3 downto 0);
    signal s3_lcd_data_low : std_logic_vector(2 downto 0) := c_LCD_REG_DATA_RESET;
    signal s3_lcd_data_high : std_logic_vector(2 downto 0) := c_LCD_REG_DATA_RESET;
    signal s_contrast : boolean := false;                                               -- Result of PWM process calculation
    signal s_backlight : boolean := false;
    signal s_bank1 : std_logic;                                                         -- Intermediate signal for controlling pout_xbox_a19 on flash chip. Will either be controlled by SW1 or OS.
    signal s_bank2 : std_logic;                                                         -- Intermediate signal for controlling A18 on flash chip. Will either be controlled by SW2 or OS.
    signal s_bank2_interm : std_logic;
    signal s_os_bnkctrl : std_logic := c_FALSE_STD;                                     -- Explicitely defined for a reason.
    signal s2_os_ctrl_bank_select : std_logic_vector(1 downto 0);                       -- OS desired bank switch state.
    signal s_os_disable : std_logic := c_FALSE_STD;                                     -- Flag raised by OS to disable modchip and boot from onboard Bios. Force complete mute until power cycle.
    signal s_temp_tsop_drv : std_logic;                                                  -- Flag raised by OS to tell modchip to control TSOP banks
    signal s_xodus_reg_base : std_logic;                                                -- Signal to identify LPC I/O) command standard to Xodus mods.
    signal s_temp_mediaboard_spoof : boolean;  
    signal s_mediaboard_spoof : boolean;                                                -- Gated to allow higher speeds. 
    signal s_mediaboard_f_nibble : boolean;
    signal s_d0_os_ctrl : std_logic := c_TRUE_STD;                                      -- Signal to toggle D0 from a LPC I/0 write command. Does not mute the modchip.
    signal s_a15_os_ctrl : std_logic := c_FALSE_STD;                                    -- Internal signal that maps to pout_xbox_a15 output IO.
    signal s_temp_tsop_bank_ctrl : std_logic := c_FALSE_STD;
    signal s_temp_tsop_drv_en : std_logic := c_FALSE_STD;
    signal s_xodus_mode : std_logic;
    signal s_enable_5v : std_logic := '0';
    signal s4_gpo : std_logic_vector(3 downto 0) := c_GPO_RESET;
    signal s_a19_ctrl : std_logic := c_FALSE_STD;
    
begin

--***+ direct signals
    pout_xbox_a19control <= s_a19_ctrl;
    s_a19_ctrl <= NOT s_temp_tsop_drv;  -- Because 74LVC125 requires a logic low signal to drive its buffer output.


    -- 256KB bank switch logic. Only upper 512KB bank is splitted into 2 256KB banks. Flash layout is as follow:
    -- 512KB(bank0) + 256KB(bank1) + 256KB(bank2) = 1MB.
    s_bank2_interm <= pin_manual_bank2 when pin_manual_bank1 = '1' and s_os_bnkctrl = c_FALSE_STD else pinout4_xbox_lad(2);
    s_bank2 <= s_bank2_interm when s_os_bnkctrl = c_FALSE_STD or s2_os_ctrl_bank_select(1) = '0'  else s2_os_ctrl_bank_select(0);
    s_bank1 <= pin_manual_bank1 when s_os_bnkctrl = c_FALSE_STD else s2_os_ctrl_bank_select(1);

    -- LCD contrast and backlight.
    pout_lcd_contrast <= '1' when s_contrast = true else '0';
    pout_lcd_backlight <= '1' when s_backlight = true else '0';

    p6out_lcd_data <= s3_lcd_data_high & s3_lcd_data_low;

    -- pout_xbox_a15 desired state mapped to output pin here.
    pout_xbox_a15 <= NOT s_a15_os_ctrl;

    pout_enable_5v <= s_enable_5v;
    p4out_gpo<= s4_gpo;

    -- Recreate LFRAME for Flash chip. Async. 
    s_lframe <= '0' when s_os_disable = c_FALSE_STD and pinout4_xbox_lad= c_LAD_START_PATTERN and s_lpc_fsm_state = LPC_FSM_WAIT_START else '1'; -- Stays at '1' when modchip is disabled. LPC flash chip will then be waiting for LFRAME to go down to start its cycle the whole time the Xbox is ON. No read from LPC then.
    pout_xbox_lframe <= s_lframe;    -- Maps to LFRAME signal on Xbox 1.6 motherboard.
    pout_flash_lframe <= s_lframe;   -- Maps to on board flash chip LFRAME signal.

    -- In both case below, replace '0' with 'Z' in case you decide to drive Xbox LFRAME/D0 signals with CPLD IO directly. A MOSFET is preferred to offer a strong signal drive.
    -- IO pin is used as VSS for LED. Do not exceed 8ma current. LED will be ON if flash read/write cycle as been detected.
    pout_n_onboard_led <= '1' when s_os_disable = c_TRUE_STD or s_d0_os_ctrl = c_FALSE_STD or s_temp_tsop_drv = c_TRUE_STD or pin_xbox_n_lrst = c_RST_ASSERTED else '0';

--***+ processes
    -- Process that cycle through all the steps of LPC RW operations. 
    processLpc : process(pin_xbox_lclk) -- 33MHz
    begin
        if rising_edge(pin_xbox_lclk) then
            if pin_xbox_n_lrst = c_RST_ASSERTED then -- Still too early in boot sequence. We must wait for RST to go high.
                s_lpc_fsm_state <= LPC_FSM_WAIT_START;   
                if s_d0_os_ctrl = c_TRUE_STD and (s_temp_tsop_drv = c_FALSE_STD or s_xodus_reg_base = c_FALSE_STD) then -- Only tie D0 to ground if not explicitly denied from OS.
                    pout_xbox_d0 <= '0';    -- Put D0 to ground.
                    if s_temp_tsop_drv = c_FALSE_STD then
                        s_xodus_mode <= c_TRUE_STD;
                    else
                        s_xodus_mode <= c_FALSE_STD;
                    end if;
                else
                    s_xodus_mode <= c_FALSE_STD;
               end if;      
            else -- There we go!
                if s_fsm_counter < c_FSM_ADDR_SEQ_NIBBLE7 then
                    s_fsm_counter <= s_fsm_counter + 1;
                else
                    s_fsm_counter <= c_FSM_COUNT_RESET;
                end if;
                case s_lpc_fsm_state is
                    when LPC_FSM_WAIT_START =>  -- 0000 read, occurs with LFRAME output asserted
                        s_io_cyc <= false;
                        if pinout4_xbox_lad = c_LAD_START_PATTERN and s_os_disable = c_FALSE_STD then -- its a start. Won't move from there if s_os_disable = '1'.
                            s_lpc_fsm_state <= LPC_FSM_GET_CYC;
                        end if;                         
                    when LPC_FSM_GET_CYC => -- next nibble is CYCTYPE
                        pout_xbox_d0 <= '1';    -- No need to hold D0 to ground now, we're already booting from LPC. 
                        if pinout4_xbox_lad(3 downto 2) = c_CYC_MEM_PREFIX then -- memory read or write
                            s_fsm_counter <= c_FSM_COUNT_RESET;    -- Reset counter for address decode.
                            s_lpc_fsm_state <= LPC_FSM_GET_ADDR;

                        elsif pinout4_xbox_lad(3 downto 2) = c_CYC_IO_PREFIX then
                            s_fsm_counter <= c_FSM_COUNT_IO_START_OFFSET;    -- Only 4 address nibbles are required in this case. IO write only requires 13 cycles.
                            s_io_cyc <= true;   -- Flag to guide state machine below into IO operations
                            s_lpc_fsm_state <= LPC_FSM_GET_ADDR;    -- LPC cycle goes on like normal.                    
                        else
                            s_lpc_fsm_state <= LPC_FSM_WAIT_START; -- sit out any unsupported cycle until the next start. This section could be expanded to allow other LPC message to go through
                        end if;
                        s_lad_dir <= pinout4_xbox_lad(1);   -- '0' is for read.
                            
                    when LPC_FSM_GET_ADDR => -- 8 nibbles of address, most significant nibble first
                        case s_fsm_counter is
                            when c_FSM_ADDR_SEQ_NIBBLE0 | c_FSM_ADDR_SEQ_NIBBLE1 =>  -- 2 first nibbles of a memory cycle must be "0xF".
                                if pinout4_xbox_lad /= c_LAD_ADDR_PATTERN1  then
                                s_lpc_fsm_state <= LPC_FSM_WAIT_START; -- sit out any unsupported cycle until the next start.
                                -- Again, this section could be expand in the event a program would want to access something else than BIOS flash.
                                end if; 
                            when c_FSM_ADDR_SEQ_NIBBLE4 =>
                                if s_io_cyc = true and pinout4_xbox_lad /= c_LAD_IOREG_PATTERN1 and pinout4_xbox_lad /= c_LAD_XODUS_PATTERN1  then -- IO cycle: first nibble must be "0xF" or "0x0"
                                        if pinout4_xbox_lad = c_LAD_MBOARD_PATTERN1 then -- 0x40** is also permitted for MediaBoard Spoof.
                                            s_temp_mediaboard_spoof <= true;
                                            s_xodus_reg_base <= c_FALSE_STD;
                                        else
                                            s_temp_mediaboard_spoof <= false;
                                            s_io_cyc <= false; -- Kick out of IO cycle state machine's branch
                                        end if;
                                else
                                    s_xodus_reg_base <= NOT pinout4_xbox_lad(3);
                                    s_temp_mediaboard_spoof <= false;
                                end if;
                            when c_FSM_ADDR_SEQ_NIBBLE5 =>
                                if s_io_cyc = true and pinout4_xbox_lad /= c_LAD_IOREG_PATTERN2 and (pinout4_xbox_lad /= c_LAD_XODUS_PATTERN2 or (s_xodus_reg_base = c_FALSE_STD and s_temp_mediaboard_spoof = false)) then     
                                    s_io_cyc <= false; -- Kick out of IO cycle state machine's branch
                                end if;
                            when c_FSM_ADDR_SEQ_NIBBLE6 =>
                                s_mediaboard_spoof <= s_temp_mediaboard_spoof; -- At this point, it is already decided if we want to spoof access to MediaBoard or not.
                                if s_temp_mediaboard_spoof = false then
                                    if s_io_cyc = true and pinout4_xbox_lad /= c_LAD_IOREG_PATTERN3 and (pinout4_xbox_lad /= c_LAD_XODUS_PATTERN3 or s_xodus_reg_base = c_FALSE_STD) then -- IO cycle: third nibble must have 3 MSBs at "000". 
                                        s_io_cyc <= false; -- Kick out of IO cycle state machine's branch
                                    end if;
                                else
                                    if pinout4_xbox_lad = c_LAD_IOREG_RD_MEDIABOARD_ID then
                                        s_mediaboard_f_nibble <= true;
                                    else
                                        s_mediaboard_f_nibble <= false;
                                    end if;
                                end if;
                            when c_FSM_ADDR_SEQ_NIBBLE7 =>
                                if s_io_cyc = true then
                                    if s_temp_mediaboard_spoof = true and s_mediaboard_f_nibble = false  then
                                        s4_io_reg_addr <=  c_LAD_IOREG_MEDIABOARD_SPOOF_GENERIC; -- Use an undefined IOREG address to feed xbox with 0x00 as data.
                                    else
                                        s4_io_reg_addr <= pinout4_xbox_lad;
                                    end if;
                                end if;
                                s_fsm_counter <= c_FSM_COUNT_RESET;
                                s_lpc_fsm_state <= LPC_FSM_DATA;
                            when others =>
                                null;
                        end case;
                    when LPC_FSM_DATA =>
                        if s_fsm_counter >= c_FSM_DATA_SEQ_MAX_COUNT then
                            s_lpc_fsm_state <= LPC_FSM_WAIT_START;
                        end if;
                    when others =>
                        null; -- How did you get there?
                end case;                   
            end if; --pin_xbox_n_lrst
        end if; -- clock
    end process processLpc;


    -- Process that control both LAD ports s_lad_dir
    -- Logic is determined by "s_lpc_fsm_state" and "s_fsm_counter" within a specific "s_lpc_fsm_state" value.
    process(s_lpc_fsm_state, s_lad_dir, s_fsm_counter, s_io_cyc, s4_io_reg_addr, p2in_gpi, s_enable_5v, s_temp_tsop_drv, s_xodus_mode, 
    s_mediaboard_f_nibble, s_a15_os_ctrl, s2_os_ctrl_bank_select, s4_gpo, pin_manual_bank1, pin_manual_bank2, s_bank1, s_bank2, s_a19_ctrl)
    begin
            if s_lpc_fsm_state = LPC_FSM_DATA and s_lad_dir = c_CYC_DIRECTION_READ and s_fsm_counter >= c_FSM_DATA_SEQ_TARA2_READ and s_fsm_counter <= c_FSM_DATA_SEQ_MAX_COUNT then -- Sequences that reverse data flow. From LPC Flash to Xbox, during read operation.
                    pinout4_flash_lad <= c_LAD_INPUT_PATTERN;
                    if s_fsm_counter = c_FSM_DATA_SEQ_SYNC_READ then
                        pinout4_xbox_lad <= c_LAD_PATTERN_SYNC; -- SYNC. Must be hard coded for IO read operations so why not use it for memory ops too.
                    else
                        if s_io_cyc = true and s_fsm_counter = c_FSM_DATA_SEQ_DATA1_READ then -- Data low nibble
                            case s4_io_reg_addr is
                                when c_LAD_IOREG_RD_DEV_ID =>
                                    if s_mediaboard_f_nibble = false then
                                        pinout4_xbox_lad <= c_DEV_ID_LOW_NIBBLE;
                                    else
                                        pinout4_xbox_lad <= c_MEDIABOARD_SPOOF_ID_LOW_NIBBLE;
                                    end if;
                                when c_LAD_IOREG_RD_MEDIABOARD_RAM =>
                                        pinout4_xbox_lad <= c_MEDIABOARD_SPOOF_RAM_SIZE;
                                when c_LAD_IOREG_RD_IO =>
                                    pinout4_xbox_lad <= p2in_gpi & s_temp_tsop_drv & s_enable_5v;
                                when c_LAD_IOREG_RD_XODUSID =>
                                    pinout4_xbox_lad <= "10" & NOT s_a15_os_ctrl & '0'; -- Spoof Chameleon modchip. Normally only maps to addr 0x00FE.
                                when c_LAD_IOREG_RD_STATUS =>
                                    -- Chameleon mode spoof
                                    -- Mode1(0x0) = Split TSOP
                                    -- Mode2(0x8) = Full TSOP
                                    -- Mode3(0x4) = 
                                    -- Mode4(0xC) = on board flash bank
                                    pinout4_xbox_lad <= NOT s_temp_tsop_drv & s_xodus_mode & s_a15_os_ctrl & s2_os_ctrl_bank_select(1);
                                when others =>
                                    pinout4_xbox_lad <= c_MEDIABOARD_SPOOF_ID_HIGH_NIBBLE;
                            end case;
                        elsif s_io_cyc = true and s_fsm_counter = c_FSM_DATA_SEQ_DATA2_READ then -- Data high nibble
                            case s4_io_reg_addr is
                                when c_LAD_IOREG_RD_DEV_ID => 
                                    if s_mediaboard_f_nibble = false then
                                        pinout4_xbox_lad <=c_DEV_ID_HIGH_NIBBLE;
                                    else
                                        pinout4_xbox_lad <= c_MEDIABOARD_SPOOF_ID_HIGH_NIBBLE;
                                    end if;
                                when c_LAD_IOREG_RD_IO =>
                                    pinout4_xbox_lad <= s4_gpo;
                                when c_LAD_IOREG_RD_XODUSID =>
                                    -- Spoof Chameleon modchip. Normally only maps to addr 0x00FE.
                                    pinout4_xbox_lad <= pin_manual_bank1 & '0' & pin_manual_bank2 & '0';    --Don't touch to the manual bank select header port for Chameleon spoof! Should be X"A".
                                when c_LAD_IOREG_RD_STATUS =>
                                    pinout4_xbox_lad <= '0' & s2_os_ctrl_bank_select(0) & s_temp_tsop_drv & s2_os_ctrl_bank_select(1);
                                when others =>
                                    pinout4_xbox_lad <= c_MEDIABOARD_SPOOF_ID_HIGH_NIBBLE;
                            end case;                                                               
                        else
                            pinout4_xbox_lad <= pinout4_flash_lad;
                        end if;
                    end if;
                    -- The rest of the time, everybody is in high-Z with pull ups so the necessary 0xF nibbles are all there.
            elsif s_lpc_fsm_state = LPC_FSM_DATA and s_lad_dir = c_CYC_DIRECTION_WRITE and s_fsm_counter >= c_FSM_DATA_SEQ_TARA2_WRITE and s_fsm_counter <= c_FSM_DATA_SEQ_MAX_COUNT  then -- Sequence that reverse data flow. From LPC Flash to Xbox, during write operation.
                    pinout4_flash_lad <= c_LAD_INPUT_PATTERN; -- Flash chip is leading the show.
                    if s_fsm_counter = c_FSM_DATA_SEQ_SYNC_WRITE then
                        pinout4_xbox_lad <= c_LAD_PATTERN_SYNC; -- SYNC. Must be hard coded for IO write operations so why not use it for memory ops too.
                    else
                        pinout4_xbox_lad <= pinout4_flash_lad;
                    end if;
                    -- The rest of the time, everybody is in high-Z with pull ups so the necessary 0xF nibbles are all there.                        
            else    -- If not one of the condition above, it means the data flow goes from the Xbox to the LPC flash. Happens on LFRAME start, CYC decode, 8 address nibbles, TARA1, TARB2 and of course when idle.
                    pinout4_xbox_lad <= c_LAD_INPUT_PATTERN;     -- Also when s_lad_dir = '1' for DATA1 and DATA2.
                    if s_lpc_fsm_state = LPC_FSM_GET_ADDR and s_fsm_counter = c_FSM_ADDR_SEQ_NIBBLE1 then
                        pinout4_flash_lad <= c_LAD_ST49LF080A_ADDR_PATTERN1;    -- Last fixed addr bit & MSB Flash chip ID
                    elsif s_lpc_fsm_state = LPC_FSM_GET_ADDR and s_fsm_counter = c_FSM_ADDR_SEQ_NIBBLE2 then 
                        pinout4_flash_lad <= c_LAD_ST49LF080A_ADDR_PATTERN2;    -- Flash chip ID bit(2) & Memory access signal bit & 2 LSB Chip ID.
                    elsif s_lpc_fsm_state = LPC_FSM_GET_ADDR and s_fsm_counter = c_FSM_ADDR_SEQ_NIBBLE3 then 
                        pinout4_flash_lad <= s_bank1 & s_bank2 & pinout4_xbox_lad(1 downto 0);  -- Nibble MSB is controlled by switch wired on "HD" solder pad. pin_manual_bank1 has external pull up so leaving this port floating will access the 
                                                                    -- higher 512KB of flash. Grounding this port will enable the lower 512KB portion of the 1MB flash.
                                                                    -- Once OS has taken control, it has priority over physical input signals
                    else
                        pinout4_flash_lad <= pinout4_xbox_lad; -- Transfer of buffer into the flash LPC port.
                    end if;     
            end if;
    end process;
    
    
    -- IO operations decoding process.
    -- Will also send the data to auxiliary output ports(p4out_gpo, LCD, etc.)
    process(pin_xbox_lclk)
    begin
    if rising_edge(pin_xbox_lclk) then
        if s_io_cyc = true and s_mediaboard_spoof = false then -- IO operation flag raised. MediaBoard doesn't have the right to talk!
                    -- Low Data nibble
                    if s_fsm_counter = c_FSM_DATA_WRITE_LO_NIBBLE_OFFSET and s_lad_dir = c_CYC_DIRECTION_WRITE then
                        case s4_io_reg_addr is
                            when c_LAD_IOREG_WR_LCD_DATA =>
                                 if s_enable_5v = '1' then
                                    s3_lcd_data_low <= pinout4_xbox_lad(3 downto 1);    
                                else
                                    s3_lcd_data_low <=  c_LCD_REG_DATA_RESET;
                                end if;
                            when c_LAD_IOREG_WR_LCD_BACKLIGHT =>
                                s6_duty_cycle_backlight(2 downto 0) <= pinout4_xbox_lad(3 downto 1); -- Skip LSB
                            when c_LAD_IOREG_WR_LCD_CONTRAST =>
                                s6_duty_cycle_contrast(2 downto 0) <= pinout4_xbox_lad(3 downto 1); -- Skip LSB
                            when c_LAD_IOREG_WR_OUTPUTS =>
                                s_enable_5v <= pinout4_xbox_lad(0);
                            when c_LAD_IOREG_WR_CTRL =>
                                s_d0_os_ctrl <= pinout4_xbox_lad(2);
                                if s_xodus_reg_base = c_TRUE_STD then
                                    s_temp_tsop_drv_en <= pinout4_xbox_lad(0);
                                    s_temp_tsop_bank_ctrl <= pinout4_xbox_lad(1);
                                    s_a15_os_ctrl <= pinout4_xbox_lad(3);
                                else
                                    s2_os_ctrl_bank_select <= pinout4_xbox_lad(1 downto 0); -- OS want to switch active flash bank
                                    pout_xbox_a19 <= pinout4_xbox_lad(3);
                                end if;
                            when others => null;
                        end case;
                        
                    -- High Data nibble  
                    elsif s_fsm_counter = c_FSM_DATA_WRITE_HI_NIBBLE_OFFSET and s_lad_dir = c_CYC_DIRECTION_WRITE then
                        case s4_io_reg_addr is
                            when c_LAD_IOREG_WR_LCD_DATA =>
                                if s_enable_5v = '1' then
                                    s3_lcd_data_high <= pinout4_xbox_lad(2 downto 0);   
                                else
                                    s3_lcd_data_high <=  c_LCD_REG_DATA_RESET;
                                end if;
                            when c_LAD_IOREG_WR_LCD_BACKLIGHT =>
                                s6_duty_cycle_backlight(5 downto 3) <= pinout4_xbox_lad(2 downto 0); 
                            when c_LAD_IOREG_WR_LCD_CONTRAST =>     
                                s6_duty_cycle_contrast(5 downto 3) <= pinout4_xbox_lad(2 downto 0);
                            when c_LAD_IOREG_WR_OUTPUTS =>
                                if s2_os_ctrl_bank_select = c_BANK_CTRL_OS_BANK and s_d0_os_ctrl = c_TRUE_STD and s_temp_tsop_drv = c_FALSE_STD then -- While we're still in OS (OS bank selected and D0 isn't manually released).
                                    s4_gpo(3 downto 2) <= pinout4_xbox_lad(3 downto 2);
                                end if;
                                s4_gpo(1 downto 0) <= pinout4_xbox_lad(1 downto 0);  
                            when c_LAD_IOREG_WR_CTRL =>
                               s_os_disable <= pinout4_xbox_lad(1); -- OS indicated to reboot from on-board BIOS. Mute modchip until power cycle.
                               if s_xodus_reg_base = c_TRUE_STD then
                                    if pinout4_xbox_lad(2) = '1' then
                                        s_temp_tsop_drv <= s_temp_tsop_drv_en;
                                        s2_os_ctrl_bank_select(1) <= s_temp_tsop_bank_ctrl;
                                        pout_xbox_a19 <= s_temp_tsop_bank_ctrl;  
                                        s2_os_ctrl_bank_select(0) <= '0';
                                    end if;
                               else
                                    s_temp_tsop_drv <= pinout4_xbox_lad(0); -- OS controls TSOP banks. 0 of this assume no control and a full TSOP load.
                                    if pinout4_xbox_lad(3) = '1' then
                                        s_os_bnkctrl <= c_TRUE_STD; -- Until power cycle. Generates warning that such signal should be set to '1' by default blablabla...
                                    end if;
                               end if;
                            when others => null;
                        end case;
                    end if;
                end if;     --s_io_cyc
            end if;     --clk
    end process;

    
    
    -- PWM processes. Generates 2 independant signals (duty cycle-wise) of a frequency of around 260KHz.
    -- Setting the duty cycle of a signal requires a single input command and will carry on the same
    -- duty cycle until a new duty cycle value is sent from the Xbox.
    process(pin_xbox_lclk)
    begin
    if(rising_edge(pin_xbox_lclk)) then
            s6_pwm_counter <= s6_pwm_counter + 1;
    end if;
    end process;    
    
    process(pin_xbox_lclk)
    begin
    if(rising_edge(pin_xbox_lclk)) then
        if s_enable_5v = '1' then
            if s6_pwm_counter = c_PWM_COUNTER_MAX_VALUE then -- Unfortunately, this code will make that even with a 0% duty cycle, signal will be set to '1' for a single cycle.
                s_backlight <= true;
            elsif s6_duty_cycle_backlight = s6_pwm_counter then
                s_backlight <= false;
            end if;
            if s6_pwm_counter = c_PWM_COUNTER_MAX_VALUE then -- Same here. So 0% Duty cycle is actually 1/64 duty cycle (1.563%).
                s_contrast <= true; -- Just toggle pout_enable_5v if you want a real 0% applied to BL and CT on the LCD!
            elsif s6_duty_cycle_contrast = s6_pwm_counter then
                s_contrast <= false;
            end if;
        else
            s_backlight <= false;
            s_contrast <= false;
        end if;
    -- That's the best I could think of to generate 2 PWM signals with 6 bits resolution each and still make it fit.
    end if;
    end process;    

end arch_lpcmod;
